.model nmos_bsim nmos level=54
+ tox=2e-9
+ u0=0.05
+ vth0=0.45
+ k1=0.53
+ k2=0.03

VGS g 0 0
VDS d 0 50m
VBS b 0 0

M1 d g 0 b nmos_bsim W=10u L=1u

.dc VGS 0 1.2 1m
.temp 300

.control
run
plot log(abs(i(VDS)))
.endc

.end
